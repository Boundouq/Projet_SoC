`ifndef OPCODES
`define OPCODES

`define INSTR_LUI     32'b???????_?????_?????_???_?????_0110111 /* LUI */
`define INSTR_AUIPC   32'b???????_?????_?????_???_?????_0010111 /* AUIPC */
`define INSTR_JAL     32'b???????_?????_?????_???_?????_1101111 /* JAL */
`define INSTR_JALR    32'b???????_?????_?????_000_?????_1100111 /* JALR */
`define INSTR_BEQ     32'b???????_?????_?????_000_?????_1100011 /* BRANCH */
`define INSTR_BNE     32'b???????_?????_?????_001_?????_1100011
`define INSTR_BLT     32'b???????_?????_?????_100_?????_1100011
`define INSTR_BGE     32'b???????_?????_?????_101_?????_1100011
`define INSTR_BLTU    32'b???????_?????_?????_110_?????_1100011
`define INSTR_BGEU    32'b???????_?????_?????_111_?????_1100011
`define INSTR_LB      32'b???????_?????_?????_000_?????_0000011 /* LOAD */
`define INSTR_LH      32'b???????_?????_?????_001_?????_0000011 //\\
`define INSTR_LW      32'b???????_?????_?????_010_?????_0000011 //\\
`define INSTR_LBU     32'b???????_?????_?????_100_?????_0000011 //\\
`define INSTR_LHU     32'b???????_?????_?????_101_?????_0000011 //\\
`define INSTR_SB      32'b???????_?????_?????_000_?????_0100011 /* STORE */
`define INSTR_SH      32'b???????_?????_?????_001_?????_0100011 //\\
`define INSTR_SW      32'b???????_?????_?????_010_?????_0100011 //\\
`define INSTR_ADDI    32'b???????_?????_?????_000_?????_0010011 /* OP-IMM */
`define INSTR_SLTI    32'b???????_?????_?????_010_?????_0010011 //\\
`define INSTR_SLTIU   32'b???????_?????_?????_011_?????_0010011 //\\
`define INSTR_XORI    32'b???????_?????_?????_100_?????_0010011 //\\
`define INSTR_ORI     32'b???????_?????_?????_110_?????_0010011 //\\
`define INSTR_ANDI    32'b???????_?????_?????_111_?????_0010011 //\\
`define INSTR_SLLI    32'b0000000_?????_?????_001_?????_0010011 //\\
`define INSTR_SRLI    32'b0000000_?????_?????_101_?????_0010011 //\\
`define INSTR_SRAI    32'b0100000_?????_?????_101_?????_0010011 //\\
`define INSTR_ADD     32'b0000000_?????_?????_000_?????_0110011 /* OP */
`define INSTR_SUB     32'b0100000_?????_?????_000_?????_0110011 //\\
`define INSTR_SLL     32'b0000000_?????_?????_001_?????_0110011 //\\
`define INSTR_SLT     32'b0000000_?????_?????_010_?????_0110011 //\\
`define INSTR_SLTU    32'b0000000_?????_?????_011_?????_0110011 //\\
`define INSTR_XOR     32'b0000000_?????_?????_100_?????_0110011 //\\
`define INSTR_SRL     32'b0000000_?????_?????_101_?????_0110011 //\\
`define INSTR_SRA     32'b0100000_?????_?????_101_?????_0110011 //\\
`define INSTR_OR      32'b0000000_?????_?????_110_?????_0110011 //\\
`define INSTR_AND     32'b0000000_?????_?????_111_?????_0110011 //\\
`define INSTR_FENCE   32'b???????_?????_?????_000_?????_0001111 /* MISC-MEM */
`define INSTR_FENCE_I 32'b???????_?????_?????_001_?????_0001111
`define INSTR_ECALL   32'b0000000_00000_00000_000_00000_1110011 /* SYSTEM */
`define INSTR_EBREAK  32'b0000000_00001_00000_000_00000_1110011
`define INSTR_MRET    32'b0011000_00010_00000_000_00000_1110011
`define INSTR_WFI     32'b0001000_00101_00000_000_00000_1110011
`define INSTR_CSRRW   32'b???????_?????_?????_001_?????_1110011
`define INSTR_CSRRS   32'b???????_?????_?????_010_?????_1110011
`define INSTR_CSRRC   32'b???????_?????_?????_011_?????_1110011
`define INSTR_CSRRWI  32'b???????_?????_?????_101_?????_1110011
`define INSTR_CSRRSI  32'b???????_?????_?????_110_?????_1110011
`define INSTR_CSRRCI  32'b???????_?????_?????_111_?????_1110011

`define INSTR_NOP     32'bxxxxxxx_xxxxx_00000_xxx_00000_0010011

`define OPCODE_JAL    7'b1101111
`define OPCODE_BRANCH 7'b1100011

`endif
