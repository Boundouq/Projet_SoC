`ifndef fetch
`define fetch


module fetch(
input req,
//input stall_in,
//input flush_in,

input instr_rvalid_in,
input gnt_in,
input [31:0] instr_rdata_in,

input branch_mispredicted_in,

output reg instr_req_out,
output reg [31:0] instr_addr_out,
output reg instr_read_out,
output reg [31:0] instr_out,
output reg [31:0] pc_out
);

reg [31:0] next_pc;
wire [31:0] pc;
assign pc = branch_mispredicted_in ? 32'b0 : next_pc;


reg [31:0] branch_offset;
assign branch_offset = 1'b1;


always @ (*) begin
  if (gnt_in) begin
    instr_req_out = 1;
    instr_addr_out = pc;
  end

end

assign instr_read_out = instr_rvalid_in;


always_ff @ (posedge req) begin
  if (instr_rvalid_in)begin
    instr_out <= instr_rdata_in;
    next_pc <= pc + branch_offset;
    pc_out <= pc;

  end
end
endmodule

`endif
